module top();


endmodule