module Control(input [5:0] OpCode,
                output reg [3:0] ALUOp,
                output reg RegWr);
    //

endmodule