module DataMemory ();


endmodule